library ieee;									--Cridem les llibreries necessaries.
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity Descodificador5 is
	Port ( Habilitacio: in STD_LOGIC;
		Ent : in STD_LOGIC_VECTOR (4 downto 0);
		Sort : out STD_LOGIC_VECTOR (31 downto 0));
end Descodificador5;

architecture desc of Descodificador5 is 

begin
	process (Habilitacio,Ent)
		begin
		if Habilitacio='1' then
		case Ent is
			when "00000" => Sort <= "00000000000000000000000000000001";
			when "00001" => Sort <= "00000000000000000000000000000010";
			when "00010" => Sort <= "00000000000000000000000000000100";
			when "00011" => Sort <= "00000000000000000000000000001000";
			when "00100" => Sort <= "00000000000000000000000000010000";
			when "00101" => Sort <= "00000000000000000000000000100000";
			when "00110" => Sort <= "00000000000000000000000001000000";
			when "00111" => Sort <= "00000000000000000000000010000000";
			when "01000" => Sort <= "00000000000000000000000100000000";
			when "01001" => Sort <= "00000000000000000000001000000000";
			when "01010" => Sort <= "00000000000000000000010000000000";
			when "01011" => Sort <= "00000000000000000000100000000000";
			when "01100" => Sort <= "00000000000000000001000000000000";
			when "01101" => Sort <= "00000000000000000010000000000000";
			when "01110" => Sort <= "00000000000000000100000000000000";
			when "01111" => Sort <= "00000000000000001000000000000000";
			when "10000" => Sort <= "00000000000000010000000000000000";
			when "10001" => Sort <= "00000000000000100000000000000000";
			when "10010" => Sort <= "00000000000001000000000000000000";
			when "10011" => Sort <= "00000000000010000000000000000000";
			when "10100" => Sort <= "00000000000100000000000000000000";
			when "10101" => Sort <= "00000000001000000000000000000000";
			when "10110" => Sort <= "00000000010000000000000000000000";
			when "10111" => Sort <= "00000000100000000000000000000000";
			when "11000" => Sort <= "00000001000000000000000000000000";
			when "11001" => Sort <= "00000010000000000000000000000000";
			when "11010" => Sort <= "00000100000000000000000000000000";
			when "11011" => Sort <= "00001000000000000000000000000000";
			when "11100" => Sort <= "00010000000000000000000000000000";
			when "11101" => Sort <= "00100000000000000000000000000000";
			when "11110" => Sort <= "01000000000000000000000000000000";
			when "11111" => Sort <= "10000000000000000000000000000000";
			when others => Sort <= "--------------------------------";
		end case;

	elsif (Habilitacio='0') then	
		Sort <= x"00000000";
		end if;
	end process;
end desc;